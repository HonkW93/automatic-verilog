$header
`timescale 1ns/1ps
module $module_name
(
);
endmodule
