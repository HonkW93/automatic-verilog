    always@(*)
    begin
         
    end
