    always@(posedge clk or negedge rst)
    begin
        if(rst==1'b1)begin
             
        end
        else begin
             
        end
    end
